-- pll.vhd

-- Generated using ACDS version 19.1 670

library IEEE;
library pll_altera_iopll_191;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity pll is
	port (
		locked   : out std_logic;        --  locked.export
		outclk_0 : out std_logic;        -- outclk0.clk
		outclk_1 : out std_logic;        -- outclk1.clk
		outclk_2 : out std_logic;        -- outclk2.clk
		refclk   : in  std_logic := '0'; --  refclk.clk
		rst      : in  std_logic := '0'  --   reset.reset
	);
end entity pll;

architecture rtl of pll is
	component pll_altera_iopll_191_zrphyuq is
		port (
			rst      : in  std_logic := 'X'; -- reset
			refclk   : in  std_logic := 'X'; -- clk
			locked   : out std_logic;        -- export
			outclk_0 : out std_logic;        -- clk
			outclk_1 : out std_logic;        -- clk
			outclk_2 : out std_logic         -- clk
		);
	end component pll_altera_iopll_191_zrphyuq;

	for iopll_0 : pll_altera_iopll_191_zrphyuq
		use entity pll_altera_iopll_191.pll_altera_iopll_191_zrphyuq;
begin

	iopll_0 : component pll_altera_iopll_191_zrphyuq
		port map (
			rst      => rst,      --   reset.reset
			refclk   => refclk,   --  refclk.clk
			locked   => locked,   --  locked.export
			outclk_0 => outclk_0, -- outclk0.clk
			outclk_1 => outclk_1, -- outclk1.clk
			outclk_2 => outclk_2  -- outclk2.clk
		);

end architecture rtl; -- of pll
