----------------------------------------------------------------------------------------------------
-- Copyright (c) ReFLEX CES 1998-2016
--
-- Use of this source code through a simulator and/or a compiler tool
-- is illegal if not authorised through ReFLEX CES License agreement.
----------------------------------------------------------------------------------------------------
----------------------------------------------------------------------------------------------------
-- Author      : Fr�d�ric Lavenant (from Jean-Louis FLOQUET entity)
-- Company     : ReFLEX CES
--               2, rue du gevaudan
--               91047 LISSES
--               FRANCE
--               http://www.reflexces.com
----------------------------------------------------------------------------------------------------
-- Description :
--
--
----------------------------------------------------------------------------------------------------
-- Version      Date            Author               Description
-- 0.1          2014/01/20      FLA                  Creation
-- 0.2          2016/10/13      JDU                 Change lib_jlf to work 
----------------------------------------------------------------------------------------------------
library ieee;
use     ieee.std_logic_1164.all;
use     ieee.numeric_std.all;

library work;
use     work.pkg_std.all;
use     work.pkg_std_unsigned.all;

package pkg_lfsr is
    function GenTaps(width : nat) return Int4Array;
    function MakeLFSR(reg : in slv) return slv;
end package pkg_lfsr;

package body pkg_lfsr is
    function GenTaps(width : nat) return Int4Array is
		variable result : Int4Array; -- Result
	begin
		result := (0,0,0,0);

		-- This table is directly extracted from the work of Ward & Milteno.
		-- This VHDL implementation requires a -1 offset on each term : this is done on final result
		case width is
			when      2 => result := (   2,   1,   0,   0);
			when      3 => result := (   3,   2,   0,   0);
			when      4 => result := (   4,   3,   0,   0);
			when      5 => result := (   5,   3,   0,   0);
			when      6 => result := (   6,   5,   0,   0);
			when      7 => result := (   7,   6,   0,   0);
			when      8 => result := (   8,   6,   5,   4);
			when      9 => result := (   9,   5,   0,   0);
			when     10 => result := (  10,   7,   0,   0);
			when     11 => result := (  11,   9,   0,   0);
			when     12 => result := (  12,  11,   8,   6);
			when     13 => result := (  13,  12,  10,   9);
			when     14 => result := (  14,  13,  11,   9);
			when     15 => result := (  15,  14,   0,   0);
			when     16 => result := (  16,  14,  13,  11);
			when     17 => result := (  17,  14,   0,   0);
			when     18 => result := (  18,  11,   0,   0);
			when     19 => result := (  19,  18,  17,  14);
			when     20 => result := (  20,  17,   0,   0);
			when     21 => result := (  21,  19,   0,   0);
			when     22 => result := (  22,  21,   0,   0);
			when     23 => result := (  23,  18,   0,   0);
			when     24 => result := (  24,  23,  21,  20);
			when     25 => result := (  25,  22,   0,   0);
			when     26 => result := (  26,  25,  24,  20);
			when     27 => result := (  27,  26,  25,  22);
			when     28 => result := (  28,  25,   0,   0);
			when     29 => result := (  29,  27,   0,   0);
			when     30 => result := (  30,  29,  26,  24);
			when     31 => result := (  31,  28,   0,   0);
			when     32 => result := (  32,  30,  26,  25);
			when     33 => result := (  33,  20,   0,   0);
			when     34 => result := (  34,  31,  30,  26);
			when     35 => result := (  35,  33,   0,   0);
			when     36 => result := (  36,  25,   0,   0);
			when     37 => result := (  37,  36,  33,  31);
			when     38 => result := (  38,  37,  33,  32);
			when     39 => result := (  39,  35,   0,   0);
			when     40 => result := (  40,  37,  36,  35);
			when     41 => result := (  41,  38,   0,   0);
			when     42 => result := (  42,  40,  37,  35);
			when     43 => result := (  43,  42,  38,  37);
			when     44 => result := (  44,  42,  39,  38);
			when     45 => result := (  45,  44,  42,  41);
			when     46 => result := (  46,  40,  39,  38);
			when     47 => result := (  47,  42,   0,   0);
			when     48 => result := (  48,  44,  41,  39);
			when     49 => result := (  49,  40,   0,   0);
			when     50 => result := (  50,  48,  47,  46);
			when     51 => result := (  51,  50,  48,  45);
			when     52 => result := (  52,  49,   0,   0);
			when     53 => result := (  53,  52,  51,  47);
			when     54 => result := (  54,  51,  48,  46);
			when     55 => result := (  55,  31,   0,   0);
			when     56 => result := (  56,  54,  52,  49);
			when     57 => result := (  57,  50,   0,   0);
			when     58 => result := (  58,  39,   0,   0);
			when     59 => result := (  59,  57,  55,  52);
			when     60 => result := (  60,  59,   0,   0);
			when     61 => result := (  61,  60,  59,  56);
			when     62 => result := (  62,  59,  57,  56);
			when     63 => result := (  63,  62,   0,   0);
			when     64 => result := (  64,  63,  61,  60);
			when     65 => result := (  65,  47,   0,   0);
			when     66 => result := (  66,  60,  58,  57);
			when     67 => result := (  67,  66,  65,  62);
			when     68 => result := (  68,  59,   0,   0);
			when     69 => result := (  69,  67,  64,  63);
			when     70 => result := (  70,  69,  67,  65);
			when     71 => result := (  71,  65,   0,   0);
			when     72 => result := (  72,  69,  63,  62);
			when     73 => result := (  73,  48,   0,   0);
			when     74 => result := (  74,  71,  70,  67);
			when     75 => result := (  75,  74,  72,  69);
			when     76 => result := (  76,  74,  72,  71);
			when     77 => result := (  77,  75,  72,  71);
			when     78 => result := (  78,  77,  76,  71);
			when     79 => result := (  79,  70,   0,   0);
			when     80 => result := (  80,  78,  76,  71);
			when     81 => result := (  81,  77,   0,   0);
			when     82 => result := (  82,  78,  76,  73);
			when     83 => result := (  83,  81,  79,  76);
			when     84 => result := (  84,  71,   0,   0);
			when     85 => result := (  85,  84,  83,  77);
			when     86 => result := (  86,  84,  81,  80);
			when     87 => result := (  87,  74,   0,   0);
			when     88 => result := (  88,  80,  79,  77);
			when     89 => result := (  89,  51,   0,   0);
			when     90 => result := (  90,  88,  87,  85);
			when     91 => result := (  91,  90,  86,  83);
			when     92 => result := (  92,  90,  87,  86);
			when     93 => result := (  93,  91,   0,   0);
			when     94 => result := (  94,  73,   0,   0);
			when     95 => result := (  95,  84,   0,   0);
			when     96 => result := (  96,  90,  87,  86);
			when     97 => result := (  97,  91,   0,   0);
			when     98 => result := (  98,  87,   0,   0);
			when     99 => result := (  99,  95,  94,  92);
			when    100 => result := ( 100,  63,   0,   0);
			when    101 => result := ( 101, 100,  95,  94);
			when    102 => result := ( 102,  99,  97,  96);
			when    103 => result := ( 103,  94,   0,   0);
			when    104 => result := ( 104, 103,  94,  93);
			when    105 => result := ( 105,  89,   0,   0);
			when    106 => result := ( 106,  91,   0,   0);
			when    107 => result := ( 107, 105,  99,  98);
			when    108 => result := ( 108,  77,   0,   0);
			when    109 => result := ( 109, 107, 105, 104);
			when    110 => result := ( 110, 109, 106, 104);
			when    111 => result := ( 111, 101,   0,   0);
			when    112 => result := ( 112, 108, 106, 101);
			when    113 => result := ( 113, 104,   0,   0);
			when    114 => result := ( 114, 113, 112, 103);
			when    115 => result := ( 115, 110, 108, 107);
			when    116 => result := ( 116, 114, 111, 110);
			when    117 => result := ( 117, 116, 115, 112);
			when    118 => result := ( 118,  85,   0,   0);
			when    119 => result := ( 119, 111,   0,   0);
			when    120 => result := ( 120, 118, 114, 111);
			when    121 => result := ( 121, 103,   0,   0);
			when    122 => result := ( 122, 121, 120, 116);
			when    123 => result := ( 123, 121,   0,   0);
			when    124 => result := ( 124,  87,   0,   0);
			when    125 => result := ( 125, 120, 119, 118);
			when    126 => result := ( 126, 124, 122, 119);
			when    127 => result := ( 127, 126,   0,   0);
			when    128 => result := ( 128, 127, 126, 121);
			when    129 => result := ( 129, 124,   0,   0);
			when    130 => result := ( 130, 127,   0,   0);
			when    131 => result := ( 131, 129, 128, 123);
			when    132 => result := ( 132, 103,   0,   0);
			when    133 => result := ( 133, 131, 125, 124);
			when    134 => result := ( 134,  77,   0,   0);
			when    135 => result := ( 135, 124,   0,   0);
			when    136 => result := ( 136, 134, 133, 128);
			when    137 => result := ( 137, 116,   0,   0);
			when    138 => result := ( 138, 137, 131, 130);
			when    139 => result := ( 139, 136, 134, 131);
			when    140 => result := ( 140, 111,   0,   0);
			when    141 => result := ( 141, 140, 135, 128);
			when    142 => result := ( 142, 121,   0,   0);
			when    143 => result := ( 143, 141, 140, 138);
			when    144 => result := ( 144, 142, 140, 137);
			when    145 => result := ( 145,  93,   0,   0);
			when    146 => result := ( 146, 144, 143, 141);
			when    147 => result := ( 147, 145, 143, 136);
			when    148 => result := ( 148, 121,   0,   0);
			when    149 => result := ( 149, 142, 140, 139);
			when    150 => result := ( 150,  97,   0,   0);
			when    151 => result := ( 151, 148,   0,   0);
			when    152 => result := ( 152, 150, 149, 146);
			when    153 => result := ( 153, 152,   0,   0);
			when    154 => result := ( 154, 153, 149, 145);
			when    155 => result := ( 155, 151, 150, 148);
			when    156 => result := ( 156, 153, 151, 147);
			when    157 => result := ( 157, 155, 152, 151);
			when    158 => result := ( 158, 153, 152, 150);
			when    159 => result := ( 159, 128,   0,   0);
			when    160 => result := ( 160, 158, 157, 155);
			when    161 => result := ( 161, 143,   0,   0);
			when    162 => result := ( 162, 158, 155, 154);
			when    163 => result := ( 163, 160, 157, 156);
			when    164 => result := ( 164, 159, 158, 152);
			when    165 => result := ( 165, 162, 157, 156);
			when    166 => result := ( 166, 164, 163, 156);
			when    167 => result := ( 167, 161,   0,   0);
			when    168 => result := ( 168, 162, 159, 152);
			when    169 => result := ( 169, 135,   0,   0);
			when    170 => result := ( 170, 147,   0,   0);
			when    171 => result := ( 171, 169, 166, 165);
			when    172 => result := ( 172, 165,   0,   0);
			when    173 => result := ( 173, 171, 168, 165);
			when    174 => result := ( 174, 161,   0,   0);
			when    175 => result := ( 175, 169,   0,   0);
			when    176 => result := ( 176, 167, 165, 164);
			when    177 => result := ( 177, 169,   0,   0);
			when    178 => result := ( 178,  91,   0,   0);
			when    179 => result := ( 179, 178, 177, 175);
			when    180 => result := ( 180, 173, 170, 168);
			when    181 => result := ( 181, 180, 175, 174);
			when    182 => result := ( 182, 181, 176, 174);
			when    183 => result := ( 183, 127,   0,   0);
			when    184 => result := ( 184, 177, 176, 175);
			when    185 => result := ( 185, 161,   0,   0);
			when    186 => result := ( 186, 180, 178, 177);
			when    187 => result := ( 187, 182, 181, 180);
			when    188 => result := ( 188, 186, 183, 182);
			when    189 => result := ( 189, 187, 184, 183);
			when    190 => result := ( 190, 188, 184, 177);
			when    191 => result := ( 191, 182,   0,   0);
			when    192 => result := ( 192, 190, 178, 177);
			when    193 => result := ( 193, 178,   0,   0);
			when    194 => result := ( 194, 107,   0,   0);
			when    195 => result := ( 195, 193, 192, 187);
			when    196 => result := ( 196, 194, 187, 185);
			when    197 => result := ( 197, 195, 193, 188);
			when    198 => result := ( 198, 133,   0,   0);
			when    199 => result := ( 199, 165,   0,   0);
			when    200 => result := ( 200, 198, 197, 195);
			when    201 => result := ( 201, 187,   0,   0);
			when    202 => result := ( 202, 147,   0,   0);
			when    203 => result := ( 203, 202, 196, 195);
			when    204 => result := ( 204, 201, 200, 194);
			when    205 => result := ( 205, 203, 200, 196);
			when    206 => result := ( 206, 201, 197, 196);
			when    207 => result := ( 207, 164,   0,   0);
			when    208 => result := ( 208, 207, 205, 199);
			when    209 => result := ( 209, 203,   0,   0);
			when    210 => result := ( 210, 207, 206, 198);
			when    211 => result := ( 211, 203, 201, 200);
			when    212 => result := ( 212, 107,   0,   0);
			when    213 => result := ( 213, 211, 208, 207);
			when    214 => result := ( 214, 213, 211, 209);
			when    215 => result := ( 215, 192,   0,   0);
			when    216 => result := ( 216, 215, 213, 209);
			when    217 => result := ( 217, 172,   0,   0);
			when    218 => result := ( 218, 207,   0,   0);
			when    219 => result := ( 219, 218, 215, 211);
			when    220 => result := ( 220, 211, 210, 208);
			when    221 => result := ( 221, 219, 215, 213);
			when    222 => result := ( 222, 220, 217, 214);
			when    223 => result := ( 223, 190,   0,   0);
			when    224 => result := ( 224, 222, 217, 212);
			when    225 => result := ( 225, 193,   0,   0);
			when    226 => result := ( 226, 223, 219, 216);
			when    227 => result := ( 227, 223, 218, 217);
			when    228 => result := ( 228, 226, 217, 216);
			when    229 => result := ( 229, 228, 225, 219);
			when    230 => result := ( 230, 224, 223, 222);
			when    231 => result := ( 231, 205,   0,   0);
			when    232 => result := ( 232, 228, 223, 221);
			when    233 => result := ( 233, 159,   0,   0);
			when    234 => result := ( 234, 203,   0,   0);
			when    235 => result := ( 235, 234, 229, 226);
			when    236 => result := ( 236, 231,   0,   0);
			when    237 => result := ( 237, 236, 233, 230);
			when    238 => result := ( 238, 237, 236, 233);
			when    239 => result := ( 239, 203,   0,   0);
			when    240 => result := ( 240, 237, 235, 232);
			when    241 => result := ( 241, 171,   0,   0);
			when    242 => result := ( 242, 241, 236, 231);
			when    243 => result := ( 243, 242, 238, 235);
			when    244 => result := ( 244, 243, 240, 235);
			when    245 => result := ( 245, 244, 241, 239);
			when    246 => result := ( 246, 245, 244, 235);
			when    247 => result := ( 247, 165,   0,   0);
			when    248 => result := ( 248, 238, 234, 233);
			when    249 => result := ( 249, 163,   0,   0);
			when    250 => result := ( 250, 147,   0,   0);
			when    251 => result := ( 251, 249, 247, 244);
			when    252 => result := ( 252, 185,   0,   0);
			when    253 => result := ( 253, 252, 247, 246);
			when    254 => result := ( 254, 253, 252, 247);
			when    255 => result := ( 255, 203,   0,   0);
			when    256 => result := ( 256, 254, 251, 246);
			when    257 => result := ( 257, 245,   0,   0);
			when    258 => result := ( 258, 175,   0,   0);
			when    259 => result := ( 259, 257, 253, 249);
			when    260 => result := ( 260, 253, 252, 250);
			when    261 => result := ( 261, 257, 255, 254);
			when    262 => result := ( 262, 258, 254, 253);
			when    263 => result := ( 263, 170,   0,   0);
			when    264 => result := ( 264, 263, 255, 254);
			when    265 => result := ( 265, 223,   0,   0);
			when    266 => result := ( 266, 219,   0,   0);
			when    267 => result := ( 267, 264, 261, 259);
			when    268 => result := ( 268, 243,   0,   0);
			when    269 => result := ( 269, 268, 263, 262);
			when    270 => result := ( 270, 217,   0,   0);
			when    271 => result := ( 271, 213,   0,   0);
			when    272 => result := ( 272, 270, 266, 263);
			when    273 => result := ( 273, 250,   0,   0);
			when    274 => result := ( 274, 207,   0,   0);
			when    275 => result := ( 275, 266, 265, 264);
			when    276 => result := ( 276, 275, 273, 270);
			when    277 => result := ( 277, 274, 271, 265);
			when    278 => result := ( 278, 273,   0,   0);
			when    279 => result := ( 279, 274,   0,   0);
			when    280 => result := ( 280, 278, 275, 271);
			when    281 => result := ( 281, 188,   0,   0);
			when    282 => result := ( 282, 247,   0,   0);
			when    283 => result := ( 283, 278, 276, 271);
			when    284 => result := ( 284, 165,   0,   0);
			when    285 => result := ( 285, 280, 278, 275);
			when    286 => result := ( 286, 217,   0,   0);
			when    287 => result := ( 287, 216,   0,   0);
			when    288 => result := ( 288, 287, 278, 277);
			when    289 => result := ( 289, 268,   0,   0);
			when    290 => result := ( 290, 288, 287, 285);
			when    291 => result := ( 291, 286, 280, 279);
			when    292 => result := ( 292, 195,   0,   0);
			when    293 => result := ( 293, 292, 287, 282);
			when    294 => result := ( 294, 233,   0,   0);
			when    295 => result := ( 295, 247,   0,   0);
			when    296 => result := ( 296, 292, 287, 285);
			when    297 => result := ( 297, 292,   0,   0);
			when    298 => result := ( 298, 294, 290, 287);
			when    299 => result := ( 299, 295, 293, 288);
			when    300 => result := ( 300, 293,   0,   0);
			when    301 => result := ( 301, 299, 296, 292);
			when    302 => result := ( 302, 261,   0,   0);
			when    303 => result := ( 303, 297, 291, 290);
			when    304 => result := ( 304, 303, 302, 293);
			when    305 => result := ( 305, 203,   0,   0);
			when    306 => result := ( 306, 305, 303, 299);
			when    307 => result := ( 307, 305, 303, 299);
			when    308 => result := ( 308, 306, 299, 293);
			when    309 => result := ( 309, 307, 302, 299);
			when    310 => result := ( 310, 309, 305, 302);
			when    311 => result := ( 311, 308, 306, 304);
			when    312 => result := ( 312, 307, 302, 301);
			when    313 => result := ( 313, 234,   0,   0);
			when    314 => result := ( 314, 299,   0,   0);
			when    315 => result := ( 315, 314, 306, 305);
			when    316 => result := ( 316, 181,   0,   0);
			when    317 => result := ( 317, 315, 313, 310);
			when    318 => result := ( 318, 313, 312, 310);
			when    319 => result := ( 319, 283,   0,   0);
			when    320 => result := ( 320, 319, 317, 316);
			when    321 => result := ( 321, 290,   0,   0);
			when    322 => result := ( 322, 255,   0,   0);
			when    323 => result := ( 323, 322, 320, 313);
			when    324 => result := ( 324, 321, 320, 318);
			when    325 => result := ( 325, 323, 320, 315);
			when    326 => result := ( 326, 325, 323, 316);
			when    327 => result := ( 327, 293,   0,   0);
			when    328 => result := ( 328, 323, 321, 319);
			when    329 => result := ( 329, 279,   0,   0);
			when    330 => result := ( 330, 328, 323, 322);
			when    331 => result := ( 331, 329, 325, 321);
			when    332 => result := ( 332, 209,   0,   0);
			when    333 => result := ( 333, 331,   0,   0);
			when    334 => result := ( 334, 333, 330, 327);
			when    335 => result := ( 335, 333, 328, 325);
			when    336 => result := ( 336, 335, 332, 329);
			when    337 => result := ( 337, 282,   0,   0);
			when    338 => result := ( 338, 336, 335, 332);
			when    339 => result := ( 339, 332, 329, 323);
			when    340 => result := ( 340, 337, 336, 329);
			when    341 => result := ( 341, 336, 330, 327);
			when    342 => result := ( 342, 217,   0,   0);
			when    343 => result := ( 343, 268,   0,   0);
			when    344 => result := ( 344, 338, 334, 333);
			when    345 => result := ( 345, 323,   0,   0);
			when    346 => result := ( 346, 344, 339, 335);
			when    347 => result := ( 347, 344, 337, 336);
			when    348 => result := ( 348, 344, 341, 340);
			when    349 => result := ( 349, 347, 344, 343);
			when    350 => result := ( 350, 297,   0,   0);
			when    351 => result := ( 351, 317,   0,   0);
			when    352 => result := ( 352, 346, 341, 339);
			when    353 => result := ( 353, 284,   0,   0);
			when    354 => result := ( 354, 349, 341, 340);
			when    355 => result := ( 355, 354, 350, 349);
			when    356 => result := ( 356, 349, 347, 346);
			when    357 => result := ( 357, 355, 347, 346);
			when    358 => result := ( 358, 351, 350, 344);
			when    359 => result := ( 359, 291,   0,   0);
			when    360 => result := ( 360, 359, 335, 334);
			when    361 => result := ( 361, 360, 357, 354);
			when    362 => result := ( 362, 299,   0,   0);
			when    363 => result := ( 363, 362, 356, 355);
			when    364 => result := ( 364, 297,   0,   0);
			when    365 => result := ( 365, 360, 359, 356);
			when    366 => result := ( 366, 337,   0,   0);
			when    367 => result := ( 367, 346,   0,   0);
			when    368 => result := ( 368, 361, 359, 351);
			when    369 => result := ( 369, 278,   0,   0);
			when    370 => result := ( 370, 231,   0,   0);
			when    371 => result := ( 371, 369, 368, 363);
			when    372 => result := ( 372, 369, 365, 357);
			when    373 => result := ( 373, 371, 366, 365);
			when    374 => result := ( 374, 369, 368, 366);
			when    375 => result := ( 375, 359,   0,   0);
			when    376 => result := ( 376, 371, 369, 368);
			when    377 => result := ( 377, 336,   0,   0);
			when    378 => result := ( 378, 335,   0,   0);
			when    379 => result := ( 379, 375, 370, 369);
			when    380 => result := ( 380, 333,   0,   0);
			when    381 => result := ( 381, 380, 379, 376);
			when    382 => result := ( 382, 301,   0,   0);
			when    383 => result := ( 383, 293,   0,   0);
			when    384 => result := ( 384, 378, 369, 368);
			when    385 => result := ( 385, 379,   0,   0);
			when    386 => result := ( 386, 303,   0,   0);
			when    387 => result := ( 387, 385, 379, 378);
			when    388 => result := ( 388, 387, 385, 374);
			when    389 => result := ( 389, 384, 380, 379);
			when    390 => result := ( 390, 301,   0,   0);
			when    391 => result := ( 391, 363,   0,   0);
			when    392 => result := ( 392, 386, 382, 379);
			when    393 => result := ( 393, 386,   0,   0);
			when    394 => result := ( 394, 259,   0,   0);
			when    395 => result := ( 395, 390, 389, 384);
			when    396 => result := ( 396, 371,   0,   0);
			when    397 => result := ( 397, 392, 387, 385);
			when    398 => result := ( 398, 393, 392, 384);
			when    399 => result := ( 399, 313,   0,   0);
			when    400 => result := ( 400, 398, 397, 395);
			when    401 => result := ( 401, 249,   0,   0);
			when    402 => result := ( 402, 399, 398, 393);
			when    403 => result := ( 403, 398, 395, 394);
			when    404 => result := ( 404, 215,   0,   0);
			when    405 => result := ( 405, 398, 397, 388);
			when    406 => result := ( 406, 249,   0,   0);
			when    407 => result := ( 407, 336,   0,   0);
			when    408 => result := ( 408, 407, 403, 401);
			when    409 => result := ( 409, 322,   0,   0);
			when    410 => result := ( 410, 407, 406, 400);
			when    411 => result := ( 411, 408, 401, 399);
			when    412 => result := ( 412, 265,   0,   0);
			when    413 => result := ( 413, 407, 406, 403);
			when    414 => result := ( 414, 405, 401, 398);
			when    415 => result := ( 415, 313,   0,   0);
			when    416 => result := ( 416, 414, 411, 407);
			when    417 => result := ( 417, 310,   0,   0);
			when    418 => result := ( 418, 417, 415, 403);
			when    419 => result := ( 419, 415, 414, 404);
			when    420 => result := ( 420, 412, 410, 407);
			when    421 => result := ( 421, 419, 417, 416);
			when    422 => result := ( 422, 273,   0,   0);
			when    423 => result := ( 423, 398,   0,   0);
			when    424 => result := ( 424, 422, 417, 415);
			when    425 => result := ( 425, 413,   0,   0);
			when    426 => result := ( 426, 415, 414, 412);
			when    427 => result := ( 427, 422, 421, 416);
			when    428 => result := ( 428, 323,   0,   0);
			when    429 => result := ( 429, 422, 421, 419);
			when    430 => result := ( 430, 419, 417, 415);
			when    431 => result := ( 431, 311,   0,   0);
			when    432 => result := ( 432, 429, 428, 419);
			when    433 => result := ( 433, 400,   0,   0);
			when    434 => result := ( 434, 429, 423, 422);
			when    435 => result := ( 435, 430, 426, 423);
			when    436 => result := ( 436, 271,   0,   0);
			when    437 => result := ( 437, 436, 435, 431);
			when    438 => result := ( 438, 373,   0,   0);
			when    439 => result := ( 439, 390,   0,   0);
			when    440 => result := ( 440, 439, 437, 436);
			when    441 => result := ( 441, 410,   0,   0);
			when    442 => result := ( 442, 440, 437, 435);
			when    443 => result := ( 443, 442, 437, 433);
			when    444 => result := ( 444, 435, 432, 431);
			when    445 => result := ( 445, 441, 439, 438);
			when    446 => result := ( 446, 341,   0,   0);
			when    447 => result := ( 447, 374,   0,   0);
			when    448 => result := ( 448, 444, 442, 437);
			when    449 => result := ( 449, 315,   0,   0);
			when    450 => result := ( 450, 371,   0,   0);
			when    451 => result := ( 451, 450, 441, 435);
			when    452 => result := ( 452, 448, 447, 446);
			when    453 => result := ( 453, 449, 447, 438);
			when    454 => result := ( 454, 449, 445, 444);
			when    455 => result := ( 455, 417,   0,   0);
			when    456 => result := ( 456, 454, 445, 433);
			when    457 => result := ( 457, 441,   0,   0);
			when    458 => result := ( 458, 255,   0,   0);
			when    459 => result := ( 459, 457, 454, 447);
			when    460 => result := ( 460, 399,   0,   0);
			when    461 => result := ( 461, 460, 455, 454);
			when    462 => result := ( 462, 389,   0,   0);
			when    463 => result := ( 463, 370,   0,   0);
			when    464 => result := ( 464, 460, 455, 441);
			when    465 => result := ( 465, 406,   0,   0);
			when    466 => result := ( 466, 460, 455, 452);
			when    467 => result := ( 467, 466, 461, 456);
			when    468 => result := ( 468, 464, 459, 453);
			when    469 => result := ( 469, 467, 464, 460);
			when    470 => result := ( 470, 321,   0,   0);
			when    471 => result := ( 471, 470,   0,   0);
			when    472 => result := ( 472, 470, 469, 461);
			when    473 => result := ( 473, 470, 467, 465);
			when    474 => result := ( 474, 283,   0,   0);
			when    475 => result := ( 475, 471, 467, 466);
			when    476 => result := ( 476, 461,   0,   0);
			when    477 => result := ( 477, 470, 462, 461);
			when    478 => result := ( 478, 357,   0,   0);
			when    479 => result := ( 479, 375,   0,   0);
			when    480 => result := ( 480, 473, 467, 464);
			when    481 => result := ( 481, 343,   0,   0);
			when    482 => result := ( 482, 477, 476, 473);
			when    483 => result := ( 483, 479, 477, 474);
			when    484 => result := ( 484, 379,   0,   0);
			when    485 => result := ( 485, 479, 469, 468);
			when    486 => result := ( 486, 481, 478, 472);
			when    487 => result := ( 487, 393,   0,   0);
			when    488 => result := ( 488, 487, 485, 484);
			when    489 => result := ( 489, 406,   0,   0);
			when    490 => result := ( 490, 271,   0,   0);
			when    491 => result := ( 491, 488, 485, 480);
			when    492 => result := ( 492, 491, 485, 484);
			when    493 => result := ( 493, 490, 488, 483);
			when    494 => result := ( 494, 357,   0,   0);
			when    495 => result := ( 495, 419,   0,   0);
			when    496 => result := ( 496, 494, 491, 480);
			when    497 => result := ( 497, 419,   0,   0);
			when    498 => result := ( 498, 495, 489, 487);
			when    499 => result := ( 499, 494, 493, 488);
			when    500 => result := ( 500, 499, 494, 490);
			when    501 => result := ( 501, 499, 497, 496);
			when    502 => result := ( 502, 498, 497, 494);
			when    503 => result := ( 503, 500,   0,   0);
			when    504 => result := ( 504, 502, 490, 483);
			when    505 => result := ( 505, 349,   0,   0);
			when    506 => result := ( 506, 411,   0,   0);
			when    507 => result := ( 507, 504, 501, 494);
			when    508 => result := ( 508, 399,   0,   0);
			when    509 => result := ( 509, 506, 502, 501);
			when    510 => result := ( 510, 501, 500, 498);
			when    511 => result := ( 511, 501,   0,   0);
			when    512 => result := ( 512, 510, 507, 504);
			when    513 => result := ( 513, 428,   0,   0);
			when    514 => result := ( 514, 511, 509, 507);
			when    515 => result := ( 515, 511, 508, 501);
			when    516 => result := ( 516, 514, 511, 509);
			when    517 => result := ( 517, 515, 507, 505);
			when    518 => result := ( 518, 485,   0,   0);
			when    519 => result := ( 519, 440,   0,   0);
			when    520 => result := ( 520, 509, 507, 503);
			when    521 => result := ( 521, 489,   0,   0);
			when    522 => result := ( 522, 518, 509, 507);
			when    523 => result := ( 523, 521, 517, 510);
			when    524 => result := ( 524, 357,   0,   0);
			when    525 => result := ( 525, 524, 521, 519);
			when    526 => result := ( 526, 525, 521, 517);
			when    527 => result := ( 527, 480,   0,   0);
			when    528 => result := ( 528, 526, 522, 517);
			when    529 => result := ( 529, 487,   0,   0);
			when    530 => result := ( 530, 527, 523, 520);
			when    531 => result := ( 531, 529, 525, 519);
			when    532 => result := ( 532, 531,   0,   0);
			when    533 => result := ( 533, 531, 530, 529);
			when    534 => result := ( 534, 533, 529, 527);
			when    535 => result := ( 535, 533, 529, 527);
			when    536 => result := ( 536, 533, 531, 529);
			when    537 => result := ( 537, 443,   0,   0);
			when    538 => result := ( 538, 537, 536, 533);
			when    539 => result := ( 539, 535, 534, 529);
			when    540 => result := ( 540, 361,   0,   0);
			when    541 => result := ( 541, 537, 531, 528);
			when    542 => result := ( 542, 540, 539, 533);
			when    543 => result := ( 543, 527,   0,   0);
			when    544 => result := ( 544, 538, 535, 531);
			when    545 => result := ( 545, 423,   0,   0);
			when    546 => result := ( 546, 545, 544, 538);
			when    547 => result := ( 547, 543, 540, 534);
			when    548 => result := ( 548, 545, 543, 538);
			when    549 => result := ( 549, 546, 545, 533);
			when    550 => result := ( 550, 357,   0,   0);
			when    551 => result := ( 551, 416,   0,   0);
			when    552 => result := ( 552, 550, 547, 532);
			when    553 => result := ( 553, 514,   0,   0);
			when    554 => result := ( 554, 551, 546, 543);
			when    555 => result := ( 555, 551, 546, 545);
			when    556 => result := ( 556, 403,   0,   0);
			when    557 => result := ( 557, 552, 551, 550);
			when    558 => result := ( 558, 553, 549, 544);
			when    559 => result := ( 559, 525,   0,   0);
			when    560 => result := ( 560, 554, 551, 549);
			when    561 => result := ( 561, 490,   0,   0);
			when    562 => result := ( 562, 560, 558, 551);
			when    563 => result := ( 563, 561, 554, 549);
			when    564 => result := ( 564, 401,   0,   0);
			when    565 => result := ( 565, 564, 559, 554);
			when    566 => result := ( 566, 413,   0,   0);
			when    567 => result := ( 567, 424,   0,   0);
			when    568 => result := ( 568, 558, 557, 551);
			when    569 => result := ( 569, 492,   0,   0);
			when    570 => result := ( 570, 503,   0,   0);
			when    571 => result := ( 571, 569, 566, 561);
			when    572 => result := ( 572, 571, 564, 560);
			when    573 => result := ( 573, 569, 567, 563);
			when    574 => result := ( 574, 561,   0,   0);
			when    575 => result := ( 575, 429,   0,   0);
			when    576 => result := ( 576, 573, 572, 563);
			when    577 => result := ( 577, 552,   0,   0);
			when    578 => result := ( 578, 562, 556, 555);
			when    579 => result := ( 579, 572, 570, 567);
			when    580 => result := ( 580, 579, 576, 574);
			when    581 => result := ( 581, 575, 574, 568);
			when    582 => result := ( 582, 497,   0,   0);
			when    583 => result := ( 583, 453,   0,   0);
			when    584 => result := ( 584, 581, 571, 570);
			when    585 => result := ( 585, 464,   0,   0);
			when    586 => result := ( 586, 584, 581, 579);
			when    587 => result := ( 587, 586, 581, 576);
			when    588 => result := ( 588, 437,   0,   0);
			when    589 => result := ( 589, 586, 585, 579);
			when    590 => result := ( 590, 497,   0,   0);
			when    591 => result := ( 591, 587, 585, 582);
			when    592 => result := ( 592, 591, 573, 568);
			when    593 => result := ( 593, 507,   0,   0);
			when    594 => result := ( 594, 575,   0,   0);
			when    595 => result := ( 595, 594, 593, 586);
			when    596 => result := ( 596, 592, 591, 590);
			when    597 => result := ( 597, 588, 585, 583);
			when    598 => result := ( 598, 597, 592, 591);
			when    599 => result := ( 599, 569,   0,   0);
			when    600 => result := ( 600, 599, 590, 589);
			when    601 => result := ( 601, 400,   0,   0);
			when    602 => result := ( 602, 596, 594, 591);
			when    603 => result := ( 603, 600, 599, 597);
			when    604 => result := ( 604, 600, 598, 589);
			when    605 => result := ( 605, 600, 598, 595);
			when    606 => result := ( 606, 602, 599, 591);
			when    607 => result := ( 607, 502,   0,   0);
			when    608 => result := ( 608, 606, 602, 585);
			when    609 => result := ( 609, 578,   0,   0);
			when    610 => result := ( 610, 483,   0,   0);
			when    611 => result := ( 611, 609, 607, 601);
			when    612 => result := ( 612, 607, 602, 598);
			when    613 => result := ( 613, 609, 603, 594);
			when    614 => result := ( 614, 613, 612, 607);
			when    615 => result := ( 615, 404,   0,   0);
			when    616 => result := ( 616, 614, 602, 597);
			when    617 => result := ( 617, 417,   0,   0);
			when    618 => result := ( 618, 615, 604, 598);
			when    619 => result := ( 619, 614, 611, 610);
			when    620 => result := ( 620, 619, 618, 611);
			when    621 => result := ( 621, 616, 615, 609);
			when    622 => result := ( 622, 325,   0,   0);
			when    623 => result := ( 623, 555,   0,   0);
			when    624 => result := ( 624, 617, 615, 612);
			when    625 => result := ( 625, 492,   0,   0);
			when    626 => result := ( 626, 623, 621, 613);
			when    627 => result := ( 627, 622, 617, 613);
			when    628 => result := ( 628, 405,   0,   0);
			when    629 => result := ( 629, 627, 624, 623);
			when    630 => result := ( 630, 628, 626, 623);
			when    631 => result := ( 631, 324,   0,   0);
			when    632 => result := ( 632, 629, 619, 613);
			when    633 => result := ( 633, 532,   0,   0);
			when    634 => result := ( 634, 319,   0,   0);
			when    635 => result := ( 635, 631, 625, 621);
			when    636 => result := ( 636, 632, 628, 623);
			when    637 => result := ( 637, 636, 628, 623);
			when    638 => result := ( 638, 637, 633, 632);
			when    639 => result := ( 639, 623,   0,   0);
			when    640 => result := ( 640, 638, 637, 626);
			when    641 => result := ( 641, 630,   0,   0);
			when    642 => result := ( 642, 523,   0,   0);
			when    643 => result := ( 643, 641, 640, 632);
			when    644 => result := ( 644, 634, 633, 632);
			when    645 => result := ( 645, 641, 637, 634);
			when    646 => result := ( 646, 397,   0,   0);
			when    647 => result := ( 647, 642,   0,   0);
			when    648 => result := ( 648, 647, 626, 625);
			when    649 => result := ( 649, 612,   0,   0);
			when    650 => result := ( 650, 647,   0,   0);
			when    651 => result := ( 651, 646, 638, 637);
			when    652 => result := ( 652, 559,   0,   0);
			when    653 => result := ( 653, 646, 645, 643);
			when    654 => result := ( 654, 649, 643, 640);
			when    655 => result := ( 655, 567,   0,   0);
			when    656 => result := ( 656, 646, 638, 637);
			when    657 => result := ( 657, 619,   0,   0);
			when    658 => result := ( 658, 603,   0,   0);
			when    659 => result := ( 659, 657, 655, 644);
			when    660 => result := ( 660, 657, 656, 648);
			when    661 => result := ( 661, 657, 650, 649);
			when    662 => result := ( 662, 365,   0,   0);
			when    663 => result := ( 663, 406,   0,   0);
			when    664 => result := ( 664, 662, 660, 649);
			when    665 => result := ( 665, 632,   0,   0);
			when    666 => result := ( 666, 664, 659, 656);
			when    667 => result := ( 667, 664, 660, 649);
			when    668 => result := ( 668, 658, 656, 651);
			when    669 => result := ( 669, 667, 665, 664);
			when    670 => result := ( 670, 517,   0,   0);
			when    671 => result := ( 671, 656,   0,   0);
			when    672 => result := ( 672, 667, 666, 661);
			when    673 => result := ( 673, 645,   0,   0);
			when    674 => result := ( 674, 671, 665, 660);
			when    675 => result := ( 675, 674, 672, 669);
			when    676 => result := ( 676, 435,   0,   0);
			when    677 => result := ( 677, 674, 673, 669);
			when    678 => result := ( 678, 675, 673, 663);
			when    679 => result := ( 679, 613,   0,   0);
			when    680 => result := ( 680, 679, 650, 645);
			when    681 => result := ( 681, 678, 672, 670);
			when    682 => result := ( 682, 681, 679, 675);
			when    683 => result := ( 683, 682, 677, 672);
			when    684 => result := ( 684, 681, 671, 666);
			when    685 => result := ( 685, 684, 682, 681);
			when    686 => result := ( 686, 489,   0,   0);
			when    687 => result := ( 687, 674,   0,   0);
			when    688 => result := ( 688, 682, 674, 669);
			when    689 => result := ( 689, 675,   0,   0);
			when    690 => result := ( 690, 687, 683, 680);
			when    691 => result := ( 691, 689, 685, 678);
			when    692 => result := ( 692, 393,   0,   0);
			when    693 => result := ( 693, 691, 685, 678);
			when    694 => result := ( 694, 691, 681, 677);
			when    695 => result := ( 695, 483,   0,   0);
			when    696 => result := ( 696, 694, 686, 673);
			when    697 => result := ( 697, 430,   0,   0);
			when    698 => result := ( 698, 483,   0,   0);
			when    699 => result := ( 699, 698, 689, 684);
			when    700 => result := ( 700, 698, 695, 694);
			when    701 => result := ( 701, 699, 697, 685);
			when    702 => result := ( 702, 665,   0,   0);
			when    703 => result := ( 703, 702, 696, 691);
			when    704 => result := ( 704, 701, 699, 692);
			when    705 => result := ( 705, 686,   0,   0);
			when    706 => result := ( 706, 697, 695, 692);
			when    707 => result := ( 707, 702, 699, 692);
			when    708 => result := ( 708, 421,   0,   0);
			when    709 => result := ( 709, 708, 706, 705);
			when    710 => result := ( 710, 709, 696, 695);
			when    711 => result := ( 711, 619,   0,   0);
			when    712 => result := ( 712, 709, 708, 707);
			when    713 => result := ( 713, 672,   0,   0);
			when    714 => result := ( 714, 691,   0,   0);
			when    715 => result := ( 715, 714, 711, 708);
			when    716 => result := ( 716, 533,   0,   0);
			when    717 => result := ( 717, 716, 710, 701);
			when    718 => result := ( 718, 717, 716, 713);
			when    719 => result := ( 719, 569,   0,   0);
			when    720 => result := ( 720, 718, 712, 709);
			when    721 => result := ( 721, 712,   0,   0);
			when    722 => result := ( 722, 491,   0,   0);
			when    723 => result := ( 723, 717, 710, 707);
			when    724 => result := ( 724, 719, 716, 711);
			when    725 => result := ( 725, 720, 719, 716);
			when    726 => result := ( 726, 721,   0,   0);
			when    727 => result := ( 727, 547,   0,   0);
			when    728 => result := ( 728, 726, 725, 724);
			when    729 => result := ( 729, 671,   0,   0);
			when    730 => result := ( 730, 583,   0,   0);
			when    731 => result := ( 731, 729, 725, 723);
			when    732 => result := ( 732, 729, 728, 725);
			when    733 => result := ( 733, 731, 726, 725);
			when    734 => result := ( 734, 724, 721, 720);
			when    735 => result := ( 735, 691,   0,   0);
			when    736 => result := ( 736, 730, 728, 723);
			when    737 => result := ( 737, 732,   0,   0);
			when    738 => result := ( 738, 391,   0,   0);
			when    739 => result := ( 739, 731, 723, 721);
			when    740 => result := ( 740, 587,   0,   0);
			when    741 => result := ( 741, 738, 733, 732);
			when    742 => result := ( 742, 741, 738, 730);
			when    743 => result := ( 743, 653,   0,   0);
			when    744 => result := ( 744, 743, 733, 731);
			when    745 => result := ( 745, 487,   0,   0);
			when    746 => result := ( 746, 395,   0,   0);
			when    747 => result := ( 747, 743, 741, 737);
			when    748 => result := ( 748, 744, 743, 733);
			when    749 => result := ( 749, 748, 743, 742);
			when    750 => result := ( 750, 746, 741, 734);
			when    751 => result := ( 751, 733,   0,   0);
			when    752 => result := ( 752, 749, 732, 731);
			when    753 => result := ( 753, 595,   0,   0);
			when    754 => result := ( 754, 735,   0,   0);
			when    755 => result := ( 755, 754, 745, 743);
			when    756 => result := ( 756, 407,   0,   0);
			when    757 => result := ( 757, 756, 751, 750);
			when    758 => result := ( 758, 757, 746, 741);
			when    759 => result := ( 759, 661,   0,   0);
			when    760 => result := ( 760, 757, 747, 734);
			when    761 => result := ( 761, 758,   0,   0);
			when    762 => result := ( 762, 679,   0,   0);
			when    763 => result := ( 763, 754, 749, 747);
			when    764 => result := ( 764, 761, 759, 758);
			when    765 => result := ( 765, 760, 755, 754);
			when    766 => result := ( 766, 757, 747, 744);
			when    767 => result := ( 767, 599,   0,   0);
			when    768 => result := ( 768, 764, 751, 749);
			when    769 => result := ( 769, 649,   0,   0);
			when    770 => result := ( 770, 768, 765, 756);
			when    771 => result := ( 771, 765, 756, 754);
			when    772 => result := ( 772, 765,   0,   0);
			when    773 => result := ( 773, 767, 765, 763);
			when    774 => result := ( 774, 589,   0,   0);
			when    775 => result := ( 775, 408,   0,   0);
			when    776 => result := ( 776, 773, 764, 759);
			when    777 => result := ( 777, 748,   0,   0);
			when    778 => result := ( 778, 403,   0,   0);
			when    779 => result := ( 779, 776, 771, 769);
			when    780 => result := ( 780, 775, 772, 764);
			when    781 => result := ( 781, 779, 765, 764);
			when    782 => result := ( 782, 453,   0,   0);
			when    783 => result := ( 783, 715,   0,   0);
			when    784 => result := ( 784, 778, 775, 771);
			when    785 => result := ( 785, 693,   0,   0);
			when    786 => result := ( 786, 782, 780, 771);
			when   1024 => result := (1024,1015,1002,1001);
			when   2048 => result := (2048,2035,2034,2029);
			when   4096 => result := (4096,4095,4081,4069);
			when others => report "[LFSR] : Unsupported WIDTH value !!" severity failure;
		end case;
		result(0) := result(0) - 1;
		result(1) := result(1) - 1;
		result(2) := result(2) - 1;
		result(3) := result(3) - 1;
		return result;
	end function GenTaps;

	function MakeLFSR(reg : in slv) return slv is
        constant    TAPS : Int4Array := GenTaps(reg'length); -- Indicate where XOR gates shall be inserted
		variable    temp : slv(reg'length-1 downto 0); -- Temporary value for output rotated vector
	begin
		-- Create vector rotation
		temp := lsb(reg) & ExcludeLSB(reg);

		-- Ignore term #3 because it's always set and doesn't generate a XOR gate
		for i in 2 downto 0 loop
			if TAPS(i)>0 then
				temp(TAPS(i)) := reg(TAPS(i)+1) xor lsb(reg);
			end if;
		end loop;
		return temp;
	end function MakeLFSR;
end package body pkg_lfsr;
