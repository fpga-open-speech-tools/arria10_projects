
module pll (
	rst,
	refclk,
	locked,
	outclk_0,
	outclk_1,
	outclk_2);	

	input		rst;
	input		refclk;
	output		locked;
	output		outclk_0;
	output		outclk_1;
	output		outclk_2;
endmodule
